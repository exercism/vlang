module main

fn proteins(strand string) ![]string {
}
