module main

fn combinations(sum int, size int, exclude []int) [][]int {
}
