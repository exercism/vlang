module main

fn can_queen_attack(white string, black string) !bool {
}
