module main

fn nth_prime(n int) !int {

}
