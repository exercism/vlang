module main

fn largest_product(digits string, span int) !int {
}
