module main

fn is_isosceles(a f64, b f64, c f64) bool {

}

fn is_equilateral(a f64, b f64, c f64) bool {

}

fn is_scalene(a f64, b f64, c f64) bool {

}