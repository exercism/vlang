module main

fn color_code(color string) int {
}

const colors = []string{}
