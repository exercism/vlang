module main

// reverse_string returns a given string in reverse order
fn reverse_string(str string) string {
	return str.reverse()
}