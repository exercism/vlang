module main

// you'll probably want this
import rand

// define the Robot struct here
struct Robot {

}

// we need a place to store all these robots!
// make sure to update all the <TYPE>s to match
// this should probably be an array or a map ;)
fn create_robot_storage() <TYPE> {
}

fn create_robot(mut robots <TYPE>) Robot {
}

fn (mut r Robot) reset(mut robots <TYPE>) {
}