module main

fn rebase(input_base int, digits []int, output_base int) ![]int {
}
