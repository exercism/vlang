module main

fn test_drinks_water() {
	assert drinks_water() == 'Norwegian'
}

fn test_owns_zebra() {
	assert owns_zebra() == 'Japanese'
}
