module main

pub fn rows(height int) [][]int {
}
