module main

pub fn square_of_sum(n u32) u32 {
}

pub fn sum_of_squares(n u32) u32 {
}

pub fn difference(n u32) u32 {
}
