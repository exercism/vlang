module main

// define the LinkedList type here
struct LinkedList {
}

// implement these methods as a minimum
pub fn (mut l LinkedList) push(value int) {
}

pub fn (mut l LinkedList) pop() int {
}

pub fn (mut l LinkedList) unshift(value int) {
}

pub fn (mut l LinkedList) shift() int {
}

pub fn (l LinkedList) count() int {
}

pub fn (mut l LinkedList) delete(value int) {
}
