module main

pub fn keep[T](array []T, predicate fn (e T) bool) []T {
}

pub fn discard[T](array []T, predicate fn (e T) bool) []T {
}
