module main

struct HighScores {
}

// build a new HighScores
pub fn HighScores.new(scores []int) HighScores {
}

pub fn (mut high_scores HighScores) scores() []int {
}

pub fn (mut high_scores HighScores) latest() int {
}

pub fn (mut high_scores HighScores) personal_best() int {
}

pub fn (mut high_scores HighScores) personal_top_three() []int {
}
