module main

fn is_paired(input string) bool {
}
