module main

fn grains_on_square(square i64) !i64 {

}

fn total_grains_on_board() i64 {
	
}