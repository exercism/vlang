module main

fn age(seconds f64, planet string) !f64 {
	// age should return an error if the planet is not one of the 8 listed
}
