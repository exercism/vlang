module main

struct LinkedList {
	// define your data structure here
}

fn new() LinkedList {

}

fn from_array(array []int) LinkedList {

}

fn (list LinkedList) is_empty() bool {

}

fn (mut list LinkedList) push(data int) {

}

fn (mut list LinkedList) pop() ?int {

}

fn (mut list LinkedList) peek() ?int {

}

fn (mut list LinkedList) to_array() []int {

}

fn (mut list LinkedList) reverse() LinkedList {

}
