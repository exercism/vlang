module main

enum Allergen as u8 {
	eggs
	peanuts
	shellfish
	strawberries
	tomatoes
	chocolate
	pollen
	cats
}

fn allergic_to(allergen Allergen, score u8) bool {
	// Please implement the `allergic_to` function
}

fn list(score u8) []Allergen {
	// Please implement the `list` function
}
