module main

fn annotate(minefield []string) []string {
}
