module main

fn truncate(phrase string) string {
}
