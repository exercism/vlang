module main

fn score(word string) int {
}
