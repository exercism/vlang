module main

pub fn is_valid(isbn_10 string) bool {
}
