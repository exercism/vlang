module main

struct Point {
	row    int
	column int
}

fn saddle_points(matrix [][]int) []Point {
}
