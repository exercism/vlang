module main

fn recite(start_verse int, end_verse int) string {
}
