module main

struct Rational {
}

// build a new Rational number
pub fn Rational.new(denominator i64, numerator i64) Rational {
}

pub fn (r Rational) abs() Rational {
}

pub fn (r Rational) add(other Rational) Rational {
}

pub fn (r Rational) div(other Rational) Rational {
}

pub fn (r Rational) exprational(n i64) Rational {
}

pub fn (r Rational) expreal(n i64) f64 {
}

pub fn (r Rational) mul(other Rational) Rational {
}

pub fn (r Rational) reduce() Rational {
}

pub fn (r Rational) sub(other Rational) Rational {
}
