module main

struct Palindrome {
	value   ?int
	factors [][]int
}

fn smallest(min int, max int) !Palindrome {
}

fn largest(min int, max int) !Palindrome {
}
