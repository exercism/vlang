module main

fn spiral_matrix(size int) [][]int {
}
