module main

fn clean(phrase string) !string {
}
