module main

enum Command as u8 {
	wink
	double_blink
	close_your_eyes
	jump
}

pub fn commands(encoded_message int) []Command {
	return []
}
