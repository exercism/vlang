module main

fn value(colors []string) int {
}
