module main

fn translate(phrase string) string {
}
