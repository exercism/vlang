module main

fn encode(integers []u32) []u8 {
}

fn decode(integers []u8) ![]u32 {
}
