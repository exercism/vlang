module main

fn label(colors []string) string {
}
