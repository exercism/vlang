module main

fn say(number i64) !string {
}
