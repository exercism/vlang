module main

fn recite(start_bottles int, take_down int) string {
}
