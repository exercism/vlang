module main

fn rows(letter rune) []string {
}
