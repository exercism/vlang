module main

fn row(str string, index int) []int {
}

fn column(str string, index int) []int {
}
