module main

fn annotate(garden []string) []string {
}
