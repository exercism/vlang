module main

fn winner(board []string) ?rune {
}
