module main

fn calculate_frequencies(texts []string) map[rune]int {
	// Please implement the `calculate_frequencies` function
}
