module main

// NOTE: there are multiple ways to accomplish this. To allow for automated
// testing, please fill out whatever type you choose for the type of roster.
// To make it easy to search, that has been replaced with <TYPE>. Good luck! :)

fn add_student(roster <TYPE>, name string, grade int) <TYPE> {
}

fn get_students_in_grade(roster <TYPE>, grade int) []string {
}

fn get_all_students(roster <TYPE>) []string {
}

// This is a helper function that should return an
// empty roster (type of your choosing)
fn create_new_roster() <TYPE> {
	return <TYPE>
}
