module main

fn count_nucleotides(strand string) !map[string]int {
}
