module main

fn transform(legacy map[int][]rune) map[rune]int {
}
