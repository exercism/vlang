module main

struct Clock {
}

fn new_clock(hour int, minute int) Clock {
}

fn (mut c Clock) add_time(minute int) {
}

fn (mut c Clock) subtract_time(minute int) {
}

fn (c Clock) string() string {
}
