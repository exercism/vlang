module main

fn total(basket []int) int {
}
