module main

fn convert(rows []string) !string {
}
