module main

fn roman(number int) string {
}
