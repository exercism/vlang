module main

fn is_pangram(phrase string) bool {

}