module main

fn recite(inputs []string) string {
}
