module main

fn date(phrase string) string {
}
