module main

struct Game {}

// build a new Game
fn Game.new() Game {
}

pub fn (mut g Game) roll(pins int) ! {
}

pub fn (g Game) score() !int {
}
