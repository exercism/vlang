module main

fn ciphertext(plaintext string) string {
}
