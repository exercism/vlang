module main

fn count_words(sentence string) map[string]int {
}
