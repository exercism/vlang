module main

fn slices(series string, slice_length int) ![]string {
}
