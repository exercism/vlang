module main

fn two_fer(name string) string {
}
