module main

fn find_fewest_coins(coins []int, target int) ![]int {
}
