module main

import arrays

enum Category as u8 {
	yacht
	ones
	twos
	threes
	fours
	fives
	sixes
	full_house
	four_of_a_kind
	little_straight
	big_straight
	choice
}

fn score(category Category, rolls []u8) int {
	// Please implement the score function
}
