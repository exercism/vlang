module main

fn plants(diagram string, student string) []string {
}
