module main

// reverse_string returns a given string in reverse order