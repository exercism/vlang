module main

fn tick(matrix [][]int) [][]int {
}
