module main

fn drinks_water() string {
	// Please implement the `drinks_water` function
}

fn owns_zebra() string {
	// Please implement the `owns_zebra` function
}
