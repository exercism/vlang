module main

pub fn tally(rows string) string {
}
