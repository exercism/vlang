module main

fn rotate(text string, shift_key int) string {
}
