module main

fn abbreviate(phrase string) string {
}
