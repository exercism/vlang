module main

fn response(hey_bob string) string {
}
