module main

struct Key {
	a int
	b int
}

fn encode(phrase string, key Key) !string {
}

fn decode(phrase string, key Key) !string {
}
