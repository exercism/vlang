module main

fn encode(phrase string) string {
}

fn decode(phrase string) string {
}
