module main

fn format(name string, number int) string {
}
