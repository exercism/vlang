module main

fn collatz(number int) !int {
}
