module main

enum Relation {
	equal
	sublist
	superlist
	unequal
}

fn compare(list_one []int, list_two []int) Relation {
}
