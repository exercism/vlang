module main

pub fn find(array []int, value int) !int {
	return 0
}
