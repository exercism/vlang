module main

fn encode(str string) string {
}

fn decode(str string) string {
}
