module main

pub fn is_armstrong_number(number i64) bool {
}
