module main

fn to_rna(dna string) string {
	// Add code here
}
