module main

fn transpose(lines []string) []string {
}
