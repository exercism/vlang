module main

type Domino = []int

fn can_chain(dominoes []Domino) bool {
}
