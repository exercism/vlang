module main

fn encode(msg string, rails int) string {
}

fn decode(msg string, rails int) string {
}
