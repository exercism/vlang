module main

fn sum(factors []int, limit int) int {
}
