module main

pub enum Number {
	perfect
	abundant
	deficient
}

// returns a `Result` type
pub fn classify(candidate int) !Number {
}
