module main

fn find_anagrams(subject string, candidates []string) []string {
}
