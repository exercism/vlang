module main

struct Item {
	weight int
	value  int
}

fn maximum_value(maximum_weight int, items []Item) int {
}
