module main

pub fn is_armstrong_number(number u32) bool {
}
