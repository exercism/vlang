module main

fn distance(a string, b string) !int {
}
