module main

fn sieve(limit int) []int {
}
