module main

fn prime_factors(n i64) []i64 {
}
