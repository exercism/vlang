module main

fn square_root(radicand u64) u64 {
}
