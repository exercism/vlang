module main

fn egg_count(number int) int {
}
