module main

fn raindrops(number int) string {
}
