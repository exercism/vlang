module main

fn answer(question string) ?int {
}
