module main

fn is_isogram(word string) bool {
}
