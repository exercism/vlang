module main

enum State as u8 {
	ongoing
	draw
	win
}

fn gamestate(board []string) !State {
}
