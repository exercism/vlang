module main

fn hello() string {
	return 'Goodbye, Mars!'
}
