module main

fn rectangles(strings []string) int {
}
