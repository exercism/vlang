module main

fn valid(value string) bool {
}
