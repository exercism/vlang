module main

fn score(x f64, y f64) int {
}
