module main

fn triplets_with_sum(n int) [][]int
