module main

fn test_hello(){
	assert hello() == "Hello, world!"
}